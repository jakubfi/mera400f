/*
	74154 4-bit to 16-bit decoder
*/

module decoder16(
	input en1_, en2_,
	input a, // LSB
	input b,
	input c,
	input d, // MSB
	output [0:15] o_
);

	always @ (*) begin
		case ({en1_, en2_, d, c, b, a})
			6'h0: o_ <= ~16'b1000000000000000;
			6'h1: o_ <= ~16'b0100000000000000;
			6'h2: o_ <= ~16'b0010000000000000;
			6'h3: o_ <= ~16'b0001000000000000;
			6'h4: o_ <= ~16'b0000100000000000;
			6'h5: o_ <= ~16'b0000010000000000;
			6'h6: o_ <= ~16'b0000001000000000;
			6'h7: o_ <= ~16'b0000000100000000;
			6'h8: o_ <= ~16'b0000000010000000;
			6'h9: o_ <= ~16'b0000000001000000;
			6'ha: o_ <= ~16'b0000000000100000;
			6'hb: o_ <= ~16'b0000000000010000;
			6'hc: o_ <= ~16'b0000000000001000;
			6'hd: o_ <= ~16'b0000000000000100;
			6'he: o_ <= ~16'b0000000000000010;
			6'hf: o_ <= ~16'b0000000000000001;
			default: o_ <= ~16'b0000000000000000;
		endcase
	end

endmodule

// vim: tabstop=2 shiftwidth=2 autoindent noexpandtab
