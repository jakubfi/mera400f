module mera400f(
	input [15:0] w,
	output [15:0] l,
	input czytrn,
	input piszrn,
	input czytrw,
	input piszrw,
	input ra, rb,
  output [0:8] r0,
  input zs, s_1, s0, carry,
  input vl, vg, exy, exx,
  input strob1,
  input ust_z, ust_v, ust_mc, ust_y, ust_x,
  input cleg,
  input w_zmvc, w_legy,
  input w8_x,
  input zero_v,
  input zer
);

endmodule

// vim: tabstop=2 shiftwidth=2 autoindent noexpandtab
